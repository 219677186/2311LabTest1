** Profile: "SCHEMATIC1-SWEEPPPP"  [ Z:\Downloads\ACSWEEP-PSpiceFiles\SCHEMATIC1\SWEEPPPP.sim ] 

** Creating circuit file "SWEEPPPP.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\adriansd\AppData\Local\Temp\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.AC DEC 11 0.1 10kHz
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
