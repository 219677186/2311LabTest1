module yMux1(z, a, b, c);
output z;
input a, b, c;
wirw notC, upper, lower;

